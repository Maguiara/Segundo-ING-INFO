

module mux4_tb;

    wire test_out, test_a, test_b;



endmodule